-- ******************************************************************************
-- 
--                   /------o
--             eccelerators
--          o------/
-- 
--  This file is an Eccelerators GmbH sample project.
-- 
--  MIT License:
--  Copyright (c) 2023 Eccelerators GmbH
-- 
--  Permission is hereby granted, free of charge, to any person obtaining a copy
--  of this software and associated documentation files (the "Software"), to deal
--  in the Software without restriction, including without limitation the rights
--  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--  copies of the Software, and to permit persons to whom the Software is
--  furnished to do so, subject to the following conditions:
-- 
--  The above copyright notice and this permission notice shall be included in all
--  copies or substantial portions of the Software.
-- 
--  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--  SOFTWARE.
-- ******************************************************************************
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Phy is
    generic(ClkPeriodIn16thNs : natural);
    port(
        Clk : in std_logic;
        Rst : in std_logic;
        SClk : out std_logic;
        MiSo : in std_logic;
        MoSi : out std_logic;
        FetchTxBytePulse : in std_logic;
        ReadyToFetchTxByte : out std_logic;
        FetchRxBytePulse : out std_logic;
        RxByteIsPending : out std_logic;
        TxByte : in std_logic_vector(7 downto 0);
        RxByte : out std_logic_vector(7 downto 0);
        CPol : in std_logic;
        CPha : in std_logic;
        SClkPeriodInNs : in std_logic_vector(9 downto 0)
    );
end entity;

architecture RTL of Phy is

    procedure incStretchCount(signal StretchCount16thNs : inout unsigned (14 downto 0); SClkPeriodNs : in unsigned (9 downto 0)) is
        variable NextStretchCount16thNs : unsigned(15 downto 0);
        variable SClkHalfPeriodNs16th : unsigned(14 downto 0);
    begin
        SClkHalfPeriodNs16th := resize(SClkPeriodNs * 8, 15);
        NextStretchCount16thNs := resize(StretchCount16thNs, 16) + to_unsigned(ClkPeriodIn16thNs, 16);
        if NextStretchCount16thNs >= SClkHalfPeriodNs16th then
            StretchCount16thNs <= to_unsigned(0, 15);
        else
            StretchCount16thNs <= resize(NextStretchCount16thNs, 15);
        end if;
    end procedure;

    signal TranceiveCount : unsigned(4 downto 0);
    signal StretchCount16thNs : unsigned(14 downto 0);
    signal TxReg : std_logic_vector(7 downto 0);
    signal RxReg : std_logic_vector(7 downto 0);
    signal SclkP : std_logic;
    signal FetchedTxByte : std_logic_vector(7 downto 0);
    signal FetchedTxByteIsPending : std_logic;

begin

    Sclk <= SclkP xor CPol;
    RxByte <= RxReg;

    prcSpiTransceive : process(Clk, Rst) is
    begin
        if Rst = '1' then
            SclkP <= '0';
            MoSi <= '0';
            ReadyToFetchTxByte <= '1';
            FetchRxBytePulse <= '0';
            TranceiveCount <= to_unsigned(30, 5);
            RxReg <= (others => '0');
            TxReg <= (others => '0');
            StretchCount16thNs <= (others => '0');
            FetchedTxByte <= (others => '0');
            FetchedTxByteIsPending <= '0';
            RxByteIsPending <= '0';
        elsif rising_edge(Clk) then
            FetchRxBytePulse <= '0'; -- default assignment
            if TranceiveCount /= 30 or StretchCount16thNs /= 0 then
                incStretchCount(StretchCount16thNs, unsigned(SClkPeriodInNs));
            end if;
            if FetchTxBytePulse then
                FetchedTxByte <= TxByte;
                FetchedTxByteIsPending <= '1';
                ReadyToFetchTxByte <= '0';
            end if;
            
            if TranceiveCount = 30 then
                if FetchedTxByteIsPending then
                    TxReg <= FetchedTxByte;
                    MoSi <= FetchedTxByte(7);
                    ReadyToFetchTxByte <= '1';
                    if Cpha = '0' then
                        TranceiveCount <= to_unsigned(31, 5);
                    else
                        TranceiveCount <= to_unsigned(31, 5);
                    end if;
                    FetchedTxByteIsPending <= '0';
                    RxByteIsPending <= '1';
                end if;
            elsif TranceiveCount = 31 then
                TranceiveCount <= to_unsigned(0, 5);
            else
                if StretchCount16thNs = 0 then
                    if Cpha then
                        case to_integer(TranceiveCount) is
                            when 0 | 2 | 4 | 6 | 8 | 10 | 12 =>
                                MoSi <= TxReg(7 - to_integer(TranceiveCount(3 downto 1)));
                                SclkP <= '1';
                                TranceiveCount <= TranceiveCount + 1;
                            when 14 =>
                                MoSi <= TxReg(7 - to_integer(TranceiveCount(3 downto 1)));
                                SclkP <= '1';
                                TranceiveCount <= TranceiveCount + 1;
                            when 1 | 3 | 5 | 7 | 9 | 11 | 13 =>
                                RxReg(7 - to_integer(TranceiveCount(3 downto 1))) <= MiSo;
                                SclkP <= '0';
                                TranceiveCount <= TranceiveCount + 1;
                            when 15 =>
                                RxReg(7 - to_integer(TranceiveCount(3 downto 1))) <= MiSo;
                                FetchRxBytePulse <= '1';
                                if FetchedTxByteIsPending then
                                    TxReg <= FetchedTxByte;
                                    ReadyToFetchTxByte <= '1';
                                    FetchedTxByteIsPending <= '0';
                                    RxByteIsPending <= '1';
                                    TranceiveCount <= to_unsigned(0, 5);
                                else
                                    RxByteIsPending <= '0';
                                    TranceiveCount <= to_unsigned(30, 5);
                                end if;
                                SclkP <= '0';
                            when others =>
                                SclkP <= '0';
                                RxByteIsPending <= '0';
                                TranceiveCount <= to_unsigned(30, 5);
                        end case;
                    else
                        case to_integer(TranceiveCount) is
                            when 0 | 2 | 4 | 6 | 8 | 10 | 12 =>
                                RxReg(7 - to_integer(TranceiveCount(3 downto 1))) <= MiSo;
                                SclkP <= '1';
                                TranceiveCount <= TranceiveCount + 1;
                            when 14 =>
                                RxReg(7 - to_integer(TranceiveCount(3 downto 1))) <= MiSo;
                                SclkP <= '1';
                                FetchRxBytePulse <= '1';
                                TranceiveCount <= TranceiveCount + 1;
                            when 1 | 3 | 5 | 7 | 9 | 11 | 13 =>
                                MoSi <= TxReg(6 - to_integer(TranceiveCount(3 downto 1)));
                                SclkP <= '0';
                                TranceiveCount <= TranceiveCount + 1;
                            when 15 =>
                                if FetchedTxByteIsPending then
                                    TxReg <= FetchedTxByte;
                                    MoSi <= FetchedTxByte(7);
                                    ReadyToFetchTxByte <= '1';
                                    if Cpha = '0' then
                                        TranceiveCount <= to_unsigned(31, 5);
                                    else
                                        TranceiveCount <= to_unsigned(31, 5);
                                    end if;
                                    FetchedTxByteIsPending <= '0';
                                    RxByteIsPending <= '1';
                                    TranceiveCount <= to_unsigned(0, 5);
                                else
                                    RxByteIsPending <= '0';
                                    TranceiveCount <= to_unsigned(30, 5);
                                end if;
                                SclkP <= '0';
                            when others =>
                                SclkP <= '0';
                                RxByteIsPending <= '0';
                                TranceiveCount <= to_unsigned(30, 5);
                        end case;
                    
                    end if;
                end if;
            end if;
        end if;
    end process;

end architecture;

-- SPI Mode CPOL CPHA     Clock Polarity in Idle State     Clock Phase Used to Sample and/or Shift the Data
--    0      0       0     Logic low                         Data sampled on rising edge and shifted out on the falling edge
--    1      0       1     Logic low                         Data sampled on the falling edge and shifted out on the rising edge
--    2      1       0     Logic high                       Data sampled on the rising edge and shifted out on the falling edge
--    3      1       1     Logic high                         Data sampled on the falling edge and shifted out on the rising edge

-- SPIMode=0, CPOL=0, CPHA=0, Data sampled on rising edge and shifted out on the falling edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15         
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .         
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .        
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________               .       :       .       :                                                                        ._______:       .                                                                                                               .___________________________________
-- ReadyToFetchTxByte                     .       |_______________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       :       .                       
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |__________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxReg                ________________n-1____|_________________________________________________________________n_____________________________________________________________|__n+1__________________________________________________________________________________________________________________________|___________n+2_____
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                             :       ._______:        _______         _______         _______         _______         _______         _______        :_______.        _______         _______         _______         _______         _______         _______         _______        :_______.        
-- SClk                 _______________________________|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |___________________ 
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)         _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                       :       .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--
--                      _______________________:_______._______:__________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- RxReg                _________________________________________________________________________________n_-1__________________________________________________________________|__n____________________________________________________________________________________________________________________________|__n+1______________________
-- 
-- 
-- ********************************************************************************************************************************************************************************************************************************************************************************************************************************
--                                                                                                                                                                                                                                                                                                                                 
-- SPIMode=2, CPOL=1, CPHA=0,  Data sampled on the rising edge and shifted out on the falling edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15       
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                             :       .       :                                                                                                       .       :                                                                                                               .       .       :        
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                                       :       .                                                                                                               .       :       :        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReadyToFetchTxByte   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________.       :_______         _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______         _______:       .___________________
-- SClk                                        :       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|        
--                                             :       .       :                                                                                                       :       .                                                                                                                       .       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______:_______._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       .       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .                                                                                                               :       .                                                                                                                       :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--                                                                                                                                                                                                                                                                                                                                 
--
-- ********************************************************************************************************************************************************************************************************************************************************************************************************************************
--
-- SPIMode=1, CPOL=0, CPHA=1, Data sampled on the falling edge and shifted out on the rising edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15         
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .         
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .        
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReadyToFetchTxByte   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                               .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |__________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                             :_______.       :_______         _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______        ._______:       . 
-- SClk                 _______________________|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |___________________________ 
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--
--
-- ****************************************************************************************************************************************************************************************************************************************************************************************************************************************
--
-- SPIMode=3, CPOL=3, CPHA=1, Data sampled on the falling edge and shifted out on the rising edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15       
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       .       :                                                                                                                       .       :        
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                                       :       .                                                                                                               .       :       :        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReadyToFetchTxByte   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________.       ._______:        _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______         _______.       :___________________________
-- SClk                                        |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       .
--                                             :       .       :                                                                                                       .       :       .                                                                                                               :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       .       :       .                                                                                                               :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________._______:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               :                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--                                                                                                                                                                                                                                                                                                                                 
