-- ******************************************************************************
-- 
--                   /------o
--             eccelerators
--          o------/
-- 
--  This file is an Eccelerators GmbH sample project.
-- 
--  MIT License:
--  Copyright (c) 2023 Eccelerators GmbH
-- 
--  Permission is hereby granted, free of charge, to any person obtaining a copy
--  of this software and associated documentation files (the "Software"), to deal
--  in the Software without restriction, including without limitation the rights
--  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--  copies of the Software, and to permit persons to whom the Software is
--  furnished to do so, subject to the following conditions:
-- 
--  The above copyright notice and this permission notice shall be included in all
--  copies or substantial portions of the Software.
-- 
--  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--  SOFTWARE.
-- ******************************************************************************
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Phy is
	generic(ClkPeriodIn16thNs : natural);
	port(
		Clk : in std_logic;
		Rst : in std_logic;
		SClk : out std_logic;
		MiSo : in std_logic;
		MoSi : out std_logic;
		DoTransceivePulse : in std_logic;
		ReleaseTxDataPulse : out std_logic;
		StoreRxDataPulse : out std_logic;
		TxByte : in std_logic_vector(7 downto 0);
		RxByte : out std_logic_vector(7 downto 0);
		CPol : in std_logic;
		CPha : in std_logic;
		SClkPeriodInNs : in std_logic_vector(9 downto 0)
	);
end entity;

architecture RTL of Phy is

	function add(count_in : in unsigned (13 downto 0); count_add : in unsigned (13 downto 0)) return unsigned is
		variable count_out : unsigned(13 downto 0);
	begin
		if resize(count_in, 15) + ClkPeriodIn16thNs < resize(count_add, 15) * 8 then
			count_out := count_in + ClkPeriodIn16thNs;
		else
			count_out := (others => '0');
		end if;
		return count_out;
	end function;

	signal TranceiveCount : unsigned(3 downto 0);
	signal StretchCount : unsigned(13 downto 0);
	signal TxShiftReg : std_logic_vector(7 downto 0);
	signal RxShiftReg : std_logic_vector(7 downto 0);

begin

	MoSi <= TxShiftReg(7);
	RxByte <= RxShiftReg;

	prcSpiTransceive : process(Clk, Rst) is
	begin
		if Rst = '1' then
			SClk <= '0';
			ReleaseTxDataPulse <= '0';
			StoreRxDataPulse <= '0';
			TranceiveCount <= to_unsigned(15, 4);
			RxShiftReg <= b"0000_0000";
			TxShiftReg <= b"0000_0000";
			StretchCount <= (others => '0');
		elsif rising_edge(Clk) then
			ReleaseTxDataPulse <= '0'; -- default assignment		
			StoreRxDataPulse <= '0'; -- default assignment	
			if DoTransceivePulse then
				TxShiftReg <= TxByte;
				if CPha then
					SClk <= not CPol;
				end if;
				StretchCount <= add(to_unsigned(0, 14), resize(unsigned(SClkPeriodInNs), 14));
				TranceiveCount <= to_unsigned(0, 4);
			else
				if TranceiveCount < to_unsigned(15, 4) then
					StretchCount <= add(StretchCount, resize(unsigned(SClkPeriodInNs), 14));
					if StretchCount = 0 then
						TranceiveCount <= TranceiveCount + 1;
						if TranceiveCount = 0 then
							if not CPha then
								SClk <= not CPol;
							end if;
							RxShiftReg(0) <= MiSo;
						elsif TranceiveCount = 1 then
							SClk <= not SClk;
							TxShiftReg(7 downto 1) <= TxShiftReg(6 downto 0);
						elsif TranceiveCount = 2 
						     or TranceiveCount = 4 
						     or TranceiveCount = 6 
						     or TranceiveCount = 8 
						     or TranceiveCount = 10 
						     or TranceiveCount = 12  then
							SClk <= not SClk;
							RxShiftReg(7 downto 1) <= RxShiftReg(6 downto 0);
							RxShiftReg(0) <= MiSo;
                        elsif TranceiveCount = 3 
                             or TranceiveCount = 5 
                             or TranceiveCount = 7 
                             or TranceiveCount = 9 
                             or TranceiveCount = 11  then					
							SClk <= not SClk;
							TxShiftReg(7 downto 1) <= TxShiftReg(6 downto 0);
						elsif TranceiveCount = 13 then
							SClk <= not SClk;
							TxShiftReg(7 downto 1) <= TxShiftReg(6 downto 0);
							ReleaseTxDataPulse <= '1';
						elsif TranceiveCount = 14 then
							SClk <= not SClk;
							RxShiftReg(7 downto 1) <= RxShiftReg(6 downto 0);
							RxShiftReg(0) <= MiSo;
							StoreRxDataPulse <= '1';
						end if;
					end if;
				else
					if StretchCount = 0 then
						SClk <= CPol;
					end if;	
				end if;
			end if;
		end if;
	end process;

end architecture;

-- SPI Mode CPOL CPHA 	Clock Polarity in Idle State 	Clock Phase Used to Sample and/or Shift the Data
--    0 	 0 	  0 	Logic low 	                    Data sampled on rising edge and shifted out on the falling edge
--    1 	 0 	  1 	Logic low 	                    Data sampled on the falling edge and shifted out on the rising edge
--    2 	 1 	  0 	Logic high                   	Data sampled on the rising edge and shifted out on the falling edge
--    3 	 1 	  1 	Logic high 	                    Data sampled on the falling edge and shifted out on the rising edge

-- SPIMode=0, CPOL=0, CPHA=0, Data sampled on rising edge and shifted out on the falling edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15         
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .         
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .        
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReleaseTxDataPulse   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |__________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                             :       ._______:        _______         _______         _______         _______         _______         _______        :_______.        _______         _______         _______         _______         _______         _______         _______        :_______.        
-- SClk                 _______________________________|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |___________________ 
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)         _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                       :       .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--
--
-- ********************************************************************************************************************************************************************************************************************************************************************************************************************************
--                                                                                                                                                                                                                                                                                                                                 
-- SPIMode=2, CPOL=1, CPHA=0,  Data sampled on the rising edge and shifted out on the falling edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15       
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                             :       .       :                                                                                                       .       :                                                                                                               .       .       :        
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                                       :       .                                                                                                               .       :       :        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReleaseTxDataPulse   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________.       :_______         _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______         _______:       .___________________
-- SClk                                        :       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|        
--                                             :       .       :                                                                                                       :       .                                                                                                                       .       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______:_______._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       .       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .                                                                                                               :       .                                                                                                                       :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--                                                                                                                                                                                                                                                                                                                                 
--
-- ********************************************************************************************************************************************************************************************************************************************************************************************************************************
--
-- SPIMode=1, CPOL=0, CPHA=1, Data sampled on the falling edge and shifted out on the rising edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15         
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .         
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .        
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReleaseTxDataPulse   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                               .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |__________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                             :_______.       :_______         _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______        ._______:       . 
-- SClk                 _______________________|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |___________________________ 
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       :       .                                                                                                                       :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               .                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--
--
-- ****************************************************************************************************************************************************************************************************************************************************************************************************************************************
--
-- SPIMode=3, CPOL=3, CPHA=1, Data sampled on the falling edge and shifted out on the rising edge
--                                        15   #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15  #   0   #   1   #   2   #   3   #   4   #   5   #   6   #   7   #   8   #   9   #  10   #   11  #   12  #   13  #   14  #   15       
--                       ______                                                                                                                                                                                                                                                                                                ____
-- nCs                         |______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________|
--    
--                      ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___     ___
-- Clk                     |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|   |___|
--                                     .       :       .       :                                                                                               .       .       :                                                                                                                       .       :        
--                                     ._______:       .       :                                                                                               .       :_______.                                                                                                               .       :       .
-- DoTransceivePulse    _______________|       |_______________________________________________________________________________________________________________________|       |___________________________________________________________________________________________________________________________________________________
--                                     .       :       .       :                                                                                                       :       .                                                                                                               .       :       :        
--                                     .       :       .       :                                                                                               ._______:       .                                                                                                               ._______:       .        
-- ReleaseTxDataPulse   _______________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________________    
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                                     .       :       .       :                                                                                               .       :_______.                                                                                                       .       .       ._______.
-- StoreRxDataPulse     _______________________________________________________________________________________________________________________________________________|       |_______________________________________________________________________________________________________________________|       |___________________
--                                     .       :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________ 
-- TxByte               _|_|_|_|_|_|_|_|__n____|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                               .       :       .                                                                                                               .       :       .        
--                      _______________________.       ._______:        _______         _______         _______         _______         _______        ._______:       ._______         _______         _______         _______         _______         _______         _______         _______.       :___________________________
-- SClk                                        |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       |_______|       .
--                                             :       .       :                                                                                                       .       :       .                                                                                                               :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________:_______._______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MoSi                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :       .       :                                                                                                       .       :       .                                                                                                               :       .        
--                      _______________________:_______._______:_______________ _______________ _______________ _______________ _______________ _______________ _______________._______ _______ _______________ _______________ _______________ _______________ _______________ _______________ _______________.___________________
-- MiSo                 _|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_|_|_|_|_
--                                             :                                                                                                                       :                                                                                                                               :       .                     
--                      _______________________:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________._______:_______._______________ _______________ _______________ _______________ _______________ _______________ _______________:_______________ ___________
-- RxShiftReg(0)        _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____bit7_______|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|___bit7________|____bit6_______|____bit5_______|____bit5_______|____bit3_______|____bit2_______|____bit1_______|____bit0_______|_|_|_|_|_|_ 
--                                             :                                                                                                                               :                                                                                                                               .
--                      _______________________:_______________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________.___________________
-- RxByte               _|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|____n__|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|_|__n+1__|_|_|_|_|_|_|_|_|_|_
--                                                                                                                                                                                                                                                                                                                                 
