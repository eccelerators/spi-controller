-- ******************************************************************************
-- 
--                   /------o
--             eccelerators
--          o------/
-- 
--  This file is an Eccelerators GmbH sample project.
-- 
--  MIT License:
--  Copyright (c) 2023 Eccelerators GmbH
-- 
--  Permission is hereby granted, free of charge, to any person obtaining a copy
--  of this software and associated documentation files (the "Software"), to deal
--  in the Software without restriction, including without limitation the rights
--  to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
--  copies of the Software, and to permit persons to whom the Software is
--  furnished to do so, subject to the following conditions:
-- 
--  The above copyright notice and this permission notice shall be included in all
--  copies or substantial portions of the Software.
-- 
--  THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
--  IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
--  FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
--  AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
--  LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
--  OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
--  SOFTWARE.
-- ******************************************************************************
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    
use work.SpiControllerIfcPackage.all;
use work.tb_pkg_bus.all;
use work.tb_pkg_signals.all;
use work.tb_pkg.all;

entity tb_top_avalon is
    generic (
        stimulus_path : string := "../tb/simstm/";
        stimulus_file : string := "TestMainAvalon.stm"
    );
end;

architecture behavioural of tb_top_avalon is

    signal simdone : std_logic := '0';
    
    signal Clk : std_logic := '0';
    signal Rst : std_logic := '1';
    signal TimeoutAck_Detected : std_logic := '0';
    signal TimeoutAck_Rec_Clear : std_logic := '0';
    
    signal executing_line : integer := 0;
    signal executing_file : text_line;
    signal marker : std_logic_vector(15 downto 0) := (others => '0');
    
    signal signals_in : t_signals_in;
    signal signals_out : t_signals_out;

    signal bus_down : t_bus_down;
    signal bus_up : t_bus_up;    
  
    signal SpiControllerIfcAvalonDown : T_SpiControllerIfcAvalonDown;
    signal SpiControllerIfcAvalonUp : T_SpiControllerIfcAvalonUp;
    signal SpiControllerIfcTrace : T_SpiControllerIfcTrace;
    
    signal SClk : std_logic;
    signal MiSo : std_logic;
    signal MoSi : std_logic;
    signal nCs : std_logic_vector(14 downto 0);
    signal WPn : std_logic;
    signal HOLDn : std_logic;
    
begin

    Rst <= transport '0' after 100 ns;
    Clk <= transport (not Clk) and (not SimDone)  after 10 ns / 2; -- 100MHz

    tb_FileIo_i : entity work.tb_simstm
        generic map (
            stimulus_path => stimulus_path,
            stimulus_file => stimulus_file          
        )
        port map (
            clk => Clk,
            rst => Rst,
            simdone => SimDone,       
            executing_line => executing_line,
            executing_file => executing_file,
            marker => marker,
            signals_in => signals_in,
            signals_out => signals_out,
            bus_down => bus_down,
            bus_up => bus_up
        );
        
    SpiControllerIfcAvalonDown.Address <= bus_down.avalonmm.address(SpiControllerIfcAvalonDown.Address'LENGTH - 1 downto 0);
    SpiControllerIfcAvalonDown.ByteEnable <= bus_down.avalonmm.byteenable;
    SpiControllerIfcAvalonDown.WriteData <= bus_down.avalonmm.writedata;
    SpiControllerIfcAvalonDown.Write <= bus_down.avalonmm.write;
    SpiControllerIfcAvalonDown.Read <= bus_down.avalonmm.read;
    
    bus_up.avalonmm.readdata <= SpiControllerIfcAvalonUp.ReadData;
    bus_up.avalonmm.waitrequest <= SpiControllerIfcAvalonUp.WaitRequest;
               
    i_SpiControllerWithAvalonBus : entity work.SpiControllerWithAvalonBus
        port map(
            Clk => Clk,
            Rst => Rst,
            SpiControllerIfcAvalonDown =>  SpiControllerIfcAvalonDown,
            SpiControllerIfcAvalonUp => SpiControllerIfcAvalonUp,
            SpiControllerIfcTrace => SpiControllerIfcTrace,
            SClk => SClk,
            MiSo => MiSo,
            MoSi => MoSi,
            nCs => nCs
        );


    WPn <= 'H';
    HOLDn <= 'H';
    MiSo <= 'H';

    -- W25Q128JVxIM: QSPI mode is off by default ( W25Q128JVxIQ: QSPI mode is on by default )
    i_W25Q128JVxIM : entity work.W25Q128JVxIM
        port map(
            CLK => SClk,
            CSn => nCs(0),
            DIO => MoSi,
            DO => MiSo,
            WPn => WPn,
            HOLDn => HOLDn
        );
  
end;